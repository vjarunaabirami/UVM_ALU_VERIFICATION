package alu_pkg;
`include "defines.sv"
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "alu_sequence_item.sv"
`include "alu_sequence.sv"
`include "alu_sequencer.sv"
`include "alu_driver.sv"
`include "alu_active_monitor.sv"
`include "alu_active_agent.sv"
`include "alu_passive_monitor.sv"
`include "alu_passive_agent.sv"
`include "alu_scoreboard.sv"
`include "alu_coverage.sv"
`include "alu_environment.sv"
`include "alu_test.sv"
endpackage
